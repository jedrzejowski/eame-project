* C:\users\adam\Pulpit\EAME.asc
R1 N002 N001 {{R1.r}}
R2 N001 N020 {{R2.r}}
R3 N020 N025 {{R3.r}}
R4 N003 N002 {{R4.r}}
R5 N019 N025 {{R5.r}}
R8 N004 N003 {{R8.r}}
R9 0 N019 {{R9.r}}
XU1 0 N001 NC_01 NC_02 N002 AD549
XU2 N027 N020 NC_03 NC_04 N025 AD549
XU3 N019 N003 NC_05 NC_06 N004 AD549
C1 N011 N004 {{C1.c}}
C2 N018 N011 {{C2.c}}
C3 NC_07 N026 {{C3.c}}
R6 N026 N004 {{R6.r}}
R7 N018 N026 {{R7.r}}
R10 N012 N011 {{R10.r}}
XU4 N018 N012 NC_08 NC_09 N012 AD549
XU5 0 N005 NC_10 NC_11 N006 AD549
XU6 0 N007 NC_12 NC_13 N008 AD549
C4 N005 N012 {{C4.c}}
R11 N006 N005 {{R11.r}}
C5 N006 N005 {{C5.c}}
C6 N021 N006 {{C6.c}}
R12 N007 N021 {{R12.r}}
C7 N008 N007 {{C7.c}}
R13 N008 N007 {{R13.r}}
R14 N015 N008 {{R14.r}}
R15 N024 N015 {{R15.r}}
R16 N017 N016 {{R16.r}}
R17 N022 N017 {{R17.r}}
C8 N024 0 {{C8.c}}
C9 N022 0 {{C9.c}}
C10 N016 N015 {{C10.c}}
C11 N013 N017 {{C11.c}}
XU8 N022 N013 NC_14 NC_15 N013 AD549
XU7 N024 N016 NC_16 NC_17 N016 AD549
R18 N023 N013 {{R18.r}}
R19 N014 N023 {{R19.r}}
R20 N010 N009 {{R20.r}}
C12 N009 N013 {{C12.c}}
C13 N014 N009 {{C13.c}}
C14 N023 0 {{C14.c}}
XU9 N014 N010 NC_18 NC_19 N010 AD549
V1 N027 0 5
.tran 5
.lib ADI1.lib
.backanno
.end
