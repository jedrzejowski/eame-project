jeden {{jeden}} eqweeq
dwa {{dwa}} eqweeq
trzy {{trzy}} eqweeq