R1 N002 IN {{R1.R}}
R2 OUT N001 IN {{R2.R}}
C1 N001 N002 100n
XU1 0 N001 V 0 Out AD549
V1 V 0 5
Vin1 IN 0 SINE(0 1 10K)
.tran 1m
.lib ADI.lib
.backanno
.end